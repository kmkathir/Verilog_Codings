//   To design Half Adder using Verilog 
//   EDA PLAYGROUND LINK : https://www.edaplayground.com/x/m4FL 

/************** Design Code *******************/
          // Gate level Description 
module half_adder(a,b,sum,carry);
  input a,b;
  output sum,carry;
  
  xor x1 (sum,a,b);
  and a1 (carry,a,b);
  
endmodule

/*******************Test Bench *********************/

module half_adder_test;
  reg a,b;
  wire sum,carry;
  
  half_adder h1 (a,b,sum,carry);
  
  initial 
    begin 
      a=0; b=0;
      #10 a=0; b=1;
      
      #10 a=1; b=0;
      
      #10 a=1; b=1;
      
     #10 $finish;
      
    end
  
      initial 
        begin
          $monitor($time,"     a=%b b=%b sum=%b carry=%b ",a,b,sum,carry);
          
        end
      
      initial
        begin
          
          $dumpfile("kathir.vcd");
          $dumpvars(0,half_adder_test);
          
        end
      
      endmodule
